module ANDGate(output wire Y,input wire A, B);

wire term0;


assign Y = A & B; //this is just a basic AND gate 


    
endmodule